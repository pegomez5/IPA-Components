`include "alu"

module UrCPU (
    input clock,
);

    reg [19:0] general_purpose_register[5:0]

endmodule
