`include "ALU.v"
`include "registers.v"

module UrCPU (
    input clock,
    input reset,
);
  
endmodule
