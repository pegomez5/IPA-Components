`include "ALU.v"
`include "registers.v"
`include "control.v"
`include "memory.v"

module UrCPU (
    input clock,
);
  
endmodule

